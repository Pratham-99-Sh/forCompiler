`timescale 10ns/1ns
`include "inv.v"
module tb;

endmodule